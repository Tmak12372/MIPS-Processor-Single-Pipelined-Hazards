LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY FORWARDING IS
	GENERIC (
		SIZE : INTEGER := 32
	);
	PORT (
        ID_EX_REGISTER_RS  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        ID_EX_REGISTER_RT  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        EX_MEM_REGWRITE    : IN STD_LOGIC;
        EX_MEM_REGISTER_RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        MEM_WB_REGISTER_RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        MEM_WB_REGWRITE    : IN STD_LOGIC;
        FORWARD_A          : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        FORWARD_B          : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END FORWARDING;

ARCHITECTURE RTL OF FORWARDING IS

BEGIN

	PROC : PROCESS (ID_EX_REGISTER_RS,ID_EX_REGISTER_RT,EX_MEM_REGWRITE,EX_MEM_REGISTER_RD,MEM_WB_REGISTER_RD,MEM_WB_REGWRITE) 
	BEGIN
		  IF (MEM_WB_REGWRITE = '1' AND (MEM_WB_REGISTER_RD /= "00000") AND NOT (EX_MEM_REGWRITE = '1' AND (EX_MEM_REGISTER_RD /= "00000") AND (EX_MEM_REGISTER_RD /= ID_EX_REGISTER_RS)) AND (MEM_WB_REGISTER_RD = ID_EX_REGISTER_RS)) THEN
				FORWARD_A <= "01";
        ELSIF (EX_MEM_REGWRITE = '1' AND (EX_MEM_REGISTER_RD /= "00000") AND (EX_MEM_REGISTER_RD = ID_EX_REGISTER_RS)) THEN
            FORWARD_A <= "10";
        ELSE
            FORWARD_A <= "00";
		END IF;

        IF (MEM_WB_REGWRITE = '1' AND (MEM_WB_REGISTER_RD /= "00000") AND NOT (EX_MEM_REGWRITE = '1' AND (EX_MEM_REGISTER_RD /= "00000") AND (EX_MEM_REGISTER_RD /= ID_EX_REGISTER_RT)) AND (MEM_WB_REGISTER_RD = ID_EX_REGISTER_RT)) THEN
            FORWARD_B <= "01";
        ELSIF (EX_MEM_REGWRITE = '1' AND (EX_MEM_REGISTER_RD /= "00000") AND (EX_MEM_REGISTER_RD = ID_EX_REGISTER_RT)) THEN
            FORWARD_B <= "10";
        ELSE
            FORWARD_B <= "00";
        END IF;
	END PROCESS;
END RTL;
