LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
LIBRARY WORK;

ENTITY REGISTERS IS
	GENERIC(
		SIZE : INTEGER := 32
	);
	PORT(
		CLK																		: IN STD_LOGIC := '0';
		REGWRITE																	: IN STD_LOGIC := '0';
		READ_REGISTER_1, READ_REGISTER_2, WRITE_REGISTER			: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		WRITE_DATA																: IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := "00000000000000000000000000000000";
		READ_DATA_1, READ_DATA_2											: OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)
	);
END REGISTERS;

ARCHITECTURE RTL OF REGISTERS IS
COMPONENT Decoder_5_32 IS 
    PORT (INPUT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
          OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END COMPONENT;

COMPONENT D_FF IS 
    PORT (CLK : IN STD_LOGIC := '0';
          EN : IN STD_LOGIC := '0';
			 IDLE : IN STD_LOGIC;
          D   : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
			 LOAD : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
          OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000"
    );
END COMPONENT;

COMPONENT MUX_32_1 IS 
    PORT (
    SEL : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    IN1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN5 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN6 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN7 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN8 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN9 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN13 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN14 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN15 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN16 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN17 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN18 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN19 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN23 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN24 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN25 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN26 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN27 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN28 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN29 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN30 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN31 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN32 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END COMPONENT;


COMPONENT REGISTER_AND IS 
    PORT (A : IN STD_LOGIC;
          B   : IN STD_LOGIC;
          F : OUT STD_LOGIC
    );
END COMPONENT;

SIGNAL DECODER_OUTPUT : STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";


TYPE MATRIX IS ARRAY(0 TO SIZE-1) OF STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
	SIGNAL Registers : MATRIX := (OTHERS => (OTHERS => '0'));								 

TYPE MATRIX1 IS ARRAY(0 TO SIZE-1) OF STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
	SIGNAL Registers1 : MATRIX := (
								 0 =>  ("00000000000000000000000000000000"),   --$zero = 0
								 1 =>  ("00000000000000000000000000000000"),  --$at = 0
								 2 =>  ("00000000000000000000000000000000"),  --$v0 = 0
								 3 =>  ("00000000000000000000000000000000"),  --$v1 = 0
								 4 =>  ("00000000000000000000000000000000"),  --$a0 = 0
								 5 =>  ("00000000000000000000000000000000"),  --$a1 = 0
								 6 =>  ("00000000000000000000000000000000"),  --$a2 = 0
								 7 =>  ("00000000000000000000000000000000"),  --$a3 = 0
								 8 =>  ("00000000000000000000000000000000"),  --$t0 = 3
								 9 =>  ("00000000000000000000000000000000"),  --$t1 = 2
								 10 => ("00000000000000000000000000000000"),  --$t2 = 2
								 11 => ("00000000000000000000000000000000"),  --$t3 = 7
								 12 => ("00000000000000000000000000000000"),  --$t4 = 0
								 13 => ("00000000000000000000000000000000"),  --$t5 = 0
								 14 => ("00000000000000000000000000000000"),  --$t6 = 0
								 15 => ("00000000000000000000000000000000"),  --$t7 = 0
								 16 => ("00000000000000000000000000000000"),  --$s0 = 12
								 17 => ("00000000000000000000000000000000"),  --$s1 = 8
								 18 => ("00000000000000000000000000000000"),  --$s2 = 8
								 19 => ("00000000000000000000000000000000"),  --$s3 = 0
								 20 => ("00000000000000000000000000000000"),  --$s4 = 0
								 21 => ("00000000000000000000000000000000"),  --$s5 = 0
								 22 => ("00000000000000000000000000000000"),  --$s6 = 0
								 23 => ("00000000000000000000000000000000"),  --$s7 = 0
								 24 => ("00000000000000000000000000000000"),  --$t8 = 0
								 25 => ("00000000000000000000000000000000"),  --$t9 = 0
								 26 => ("00000000000000000000000000000000"),  --$k0 = 0
								 27 => ("00000000000000000000000000000000"),  --$k1 = 0
								 28 => ("00000000000000000000000000000000"),  --$gp = 0
								 29 => ("00000000000000000000000000000000"),  --$sp = 0
								 30 => ("00000000000000000000000000000000"),  --$fp = 0
								 31 => ("00000000000000000000000000000000"),  --$ra = 0
								 OTHERS => (OTHERS => '0'));
								 
								 
								 
TYPE MAT IS ARRAY(0 TO SIZE-1) OF STD_LOGIC;
	SIGNAL C : MAT := (OTHERS => '0');
								





	signal IsStartup : STD_LOGIC := '1';

BEGIN
	
	process(CLK)
	begin
	  if rising_edge(CLK) then
		 IsStartup <= '0';
	  end if;
	end process;
	
    U50 : Decoder_5_32 PORT MAP (WRITE_REGISTER,DECODER_OUTPUT);

	 GEN1 : for i in 0 to 31 generate
		U51 : REGISTER_AND PORT MAP(REGWRITE,DECODER_OUTPUT(i),C(i));
	 end generate;
	 
	 GEN2 : for i in 0 to 31 generate
		U90 : D_FF PORT MAP (CLK,C(i),IsStartup,WRITE_DATA,REGISTERS1(i),REGISTERS(i));
	 end generate;
	 
    U122 : MUX_32_1 PORT MAP (READ_REGISTER_1,REGISTERS(0),REGISTERS(1),REGISTERS(2),REGISTERS(3),REGISTERS(4),REGISTERS(5),REGISTERS(6),REGISTERS(7),REGISTERS(8),REGISTERS(9),REGISTERS(10),REGISTERS(11),REGISTERS(12),REGISTERS(13),REGISTERS(14),REGISTERS(15),REGISTERS(16),REGISTERS(17),REGISTERS(18),REGISTERS(19),REGISTERS(20),REGISTERS(21),REGISTERS(22),REGISTERS(23),REGISTERS(24),REGISTERS(25),REGISTERS(26),REGISTERS(27),REGISTERS(28),REGISTERS(29),REGISTERS(30),REGISTERS(31),READ_DATA_1);
    U123 : MUX_32_1 PORT MAP (READ_REGISTER_2,REGISTERS(0),REGISTERS(1),REGISTERS(2),REGISTERS(3),REGISTERS(4),REGISTERS(5),REGISTERS(6),REGISTERS(7),REGISTERS(8),REGISTERS(9),REGISTERS(10),REGISTERS(11),REGISTERS(12),REGISTERS(13),REGISTERS(14),REGISTERS(15),REGISTERS(16),REGISTERS(17),REGISTERS(18),REGISTERS(19),REGISTERS(20),REGISTERS(21),REGISTERS(22),REGISTERS(23),REGISTERS(24),REGISTERS(25),REGISTERS(26),REGISTERS(27),REGISTERS(28),REGISTERS(29),REGISTERS(30),REGISTERS(31),READ_DATA_2);
	 
	 
	 
	 END RTL;