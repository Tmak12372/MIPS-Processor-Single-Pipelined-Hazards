LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TESTBENCH IS
END TESTBENCH;

ARCHITECTURE RTL OF TESTBENCH IS
COMPONENT MIPS_PROCESSOR IS
	GENERIC(
		SIZE : INTEGER := 32
		);
	PORT (
		CLK 			 	 : IN STD_LOGIC;
		O_REG_WRITTEN     : OUT STD_LOGIC;
		O_INSTRUCTION_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		O_RD					 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		O_RS 				 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		O_RT					 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		O_PC_OUTPUT 		 : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		O_ALU_RESULT      : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)		
		);

END COMPONENT;
	
COMPONENT REGISTERS IS
	GENERIC(
		SIZE : INTEGER := 32
	);
	PORT(
		CLK																		: IN STD_LOGIC;
		REGWRITE																	: IN STD_LOGIC;
		READ_REGISTER_1, READ_REGISTER_2, WRITE_REGISTER			: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		WRITE_DATA																: IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		READ_DATA_1, READ_DATA_2											: OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)
	);
END COMPONENT;	
	
	SIGNAL CLK_TB,STOP_BIT,REG_WRITTEN_TB : STD_LOGIC := '0';
	SIGNAL NUM_ADD_TB : STD_LOGIC_VECTOR(2 DOWNTO 0) := "100";
	SIGNAL RD_TB,RS_TB,RT_TB : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
	SIGNAL PC_OUT_TB : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL INSTRUCTION_OUT_TB,ALU_RESULT_TB : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	--SIGNAL WRITE_DATA_TB,READ_DATA_1_TB,READ_DATA_2_TB : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	
BEGIN

	UUT : MIPS_PROCESSOR PORT MAP(CLK_TB,REG_WRITTEN_TB,INSTRUCTION_OUT_TB,RD_TB,RS_TB,RT_TB,PC_OUT_TB,ALU_RESULT_TB);
	--UUT1 : REGISTERS PORT MAP(CLK_TB,REG_WRITTEN_TB,RS_TB,RT_TB,RD_TB,WRITE_DATA_TB,READ_DATA_1_TB,READ_DATA_2_TB);
	CLK_1 : PROCESS
		BEGIN
			CLK_TB <= '0'; WAIT FOR 10NS;
			CLK_TB <= '1'; WAIT FOR 10NS;
			IF (STOP_BIT = '1') THEN
				WAIT;
			END IF;
			
	END PROCESS;
	
	STIMULUS : PROCESS
	BEGIN
		
		WAIT FOR 120NS;
		STOP_BIT <= '1'; --USED FOR GOING THROUGH INSTRUCTIONS
		WAIT;
	END PROCESS;
	
END RTL;