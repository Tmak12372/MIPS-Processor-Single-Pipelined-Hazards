LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY AND_GATE IS		
	PORT (
		A : IN STD_LOGIC;
        B : IN STD_LOGIC;
		F : OUT STD_LOGIC);
END AND_GATE;

ARCHITECTURE RTL OF AND_GATE IS
BEGIN
	PROC : PROCESS (A,B) 
	BEGIN
		IF (A = '1' AND B = '1') THEN
            F <= '1';
        ELSE 
            F <= '0';
        END IF;
	END PROCESS;
END RTL;
