LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY PROGRAM_COUNTER IS
	GENERIC (
		SIZE : INTEGER := 32
		);
		
	PORT (
		CLK 		: IN STD_LOGIC;
		ADDRESS_IN  : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := (OTHERS => '0');
		ADDRESS_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := (OTHERS => '0')
		);
END PROGRAM_COUNTER;

ARCHITECTURE RTL OF PROGRAM_COUNTER IS

BEGIN

	PROC : PROCESS (CLK,ADDRESS_IN) --SYNCHRONOUS SYSTEM
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
			ADDRESS_OUT <= ADDRESS_IN; --DFF that holds our program counter 
		END IF;
	END PROCESS;
END RTL;
