LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
LIBRARY WORK;

ENTITY MIPS_PROCESSOR IS
	GENERIC(
		SIZE : INTEGER := 32; --Makes changing size easier 
		ADDR_SIZE : INTEGER := 8
		);
	PORT (
		CLK 			: IN STD_LOGIC := '0'; 
		INSTRUCTION_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		PC_INPUT 	: OUT STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		PC_OUTPUT 		: OUT STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		READ_ADDRESS : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0')
	);

END MIPS_PROCESSOR;

ARCHITECTURE RTL OF MIPS_PROCESSOR IS
	SIGNAL PC_ADDR_INPUT, PC_ADDR_OUTPUT : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL IP_TO_INST : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL IR_ADDR_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL IP_Q : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL RESET : STD_LOGIC;
BEGIN

	U1 : ENTITY WORK.PROGRAM_COUNTER PORT MAP(CLK,PC_ADDR_INPUT,PC_ADDR_OUTPUT); --Program counter 
	U2 : ENTITY WORK.ADDER PORT MAP(PC_ADDR_OUTPUT,PC_ADDR_INPUT); --Increments the Program counter
	U3 : ENTITY WORK.IP_MEMORY PORT MAP(PC_ADDR_OUTPUT(7 DOWNTO 0),CLK, x"00000000", '0',IP_Q); --Brings in instructions from a .mif file
	
	INSTRUCTION_OUT <= IP_Q; --FOR TESTBENCH
	READ_ADDRESS <= PC_ADDR_OUTPUT(7 DOWNTO 0);
	PC_INPUT <= PC_ADDR_INPUT(5 DOWNTO 0); --FOR TESTBENCH
	PC_OUTPUT <= PC_ADDR_OUTPUT(5 DOWNTO 0); --FOR TESTBENCH
END RTL;