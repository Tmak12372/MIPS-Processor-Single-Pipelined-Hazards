LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TESTBENCH IS
END TESTBENCH;

ARCHITECTURE RTL OF TESTBENCH IS
	COMPONENT MIPS_PROCESSOR IS
		GENERIC(
			SIZE : INTEGER := 32
			);
		PORT (
			CLK : IN STD_LOGIC := '0'; 
			INSTRUCTION_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			IP_OUTPUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			ADDER_OUTPUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			PC_OUTPUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			IR_ADDR_OUTPUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
			);

	END COMPONENT;
	
	
	SIGNAL CLK_TB,STOP_BIT : STD_LOGIC := '0';
	SIGNAL IP_OUT_TB,ADDER_OUT_TB,PC_OUT_TB : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL IR_ADDR_OUTPUT_TB : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL INSTRUCTION_OUT_TB : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
BEGIN
	UUT : MIPS_PROCESSOR PORT MAP(CLK_TB,INSTRUCTION_OUT_TB,IP_OUT_TB,ADDER_OUT_TB,PC_OUT_TB,IR_ADDR_OUTPUT_TB);
	CLK_1 : PROCESS
		BEGIN
			
			CLK_TB <= '1'; WAIT FOR 10NS;
			CLK_TB <= '0'; WAIT FOR 10NS;
			
			IF (STOP_BIT = '1') THEN
				WAIT;
			END IF;
			
	END PROCESS;
	
	STIMULUS : PROCESS
	BEGIN
		
		WAIT FOR 140NS;
		STOP_BIT <= '1';
		WAIT;
	END PROCESS;
	
END RTL;