LIBRARY  IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY Decoder_5_32 IS 
    PORT (INPUT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
          OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END Decoder_5_32;

ARCHITECTURE RTL OF Decoder_5_32 IS
BEGIN
    OUTPUT <= "00000000000000000000000000000001" WHEN INPUT = "00000" ELSE 
				  "00000000000000000000000000000010" WHEN INPUT = "00001" ELSE 
				  "00000000000000000000000000000100" WHEN INPUT = "00010" ELSE
				  "00000000000000000000000000001000" WHEN INPUT = "00011" ELSE
				  "00000000000000000000000000010000" WHEN INPUT = "00100" ELSE
				  "00000000000000000000000000100000" WHEN INPUT = "00101" ELSE
				  "00000000000000000000000001000000" WHEN INPUT = "00110" ELSE
				  "00000000000000000000000010000000" WHEN INPUT = "00111" ELSE
				  "00000000000000000000000100000000" WHEN INPUT = "01000" ELSE
				  "00000000000000000000001000000000" WHEN INPUT = "01001" ELSE
				  "00000000000000000000010000000000" WHEN INPUT = "01010" ELSE
				  "00000000000000000000100000000000" WHEN INPUT = "01011" ELSE
				  "00000000000000000001000000000000" WHEN INPUT = "01100" ELSE
				  "00000000000000000010000000000000" WHEN INPUT = "01101" ELSE
				  "00000000000000000100000000000000" WHEN INPUT = "01110" ELSE
				  "00000000000000001000000000000000" WHEN INPUT = "01111" ELSE
				  "00000000000000010000000000000000" WHEN INPUT = "10000" ELSE
				  "00000000000000100000000000000000" WHEN INPUT = "10001" ELSE
				  "00000000000001000000000000000000" WHEN INPUT = "10010" ELSE
				  "00000000000010000000000000000000" WHEN INPUT = "10011" ELSE
				  "00000000000100000000000000000000" WHEN INPUT = "10100" ELSE
				  "00000000001000000000000000000000" WHEN INPUT = "10101" ELSE
				  "00000000010000000000000000000000" WHEN INPUT = "10110" ELSE
				  "00000000100000000000000000000000" WHEN INPUT = "10111" ELSE
				  "00000001000000000000000000000000" WHEN INPUT = "11000" ELSE
				  "00000010000000000000000000000000" WHEN INPUT = "11001" ELSE
				  "00000100000000000000000000000000" WHEN INPUT = "11010" ELSE
				  "00001000000000000000000000000000" WHEN INPUT = "11011" ELSE
				  "00010000000000000000000000000000" WHEN INPUT = "11100" ELSE
				  "00100000000000000000000000000000" WHEN INPUT = "11101" ELSE
				  "01000000000000000000000000000000" WHEN INPUT = "11110" ELSE
				  "10000000000000000000000000000000" WHEN INPUT = "11111" ELSE
				  "00000000000000000000000000000001";
END RTL;




