LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALU IS
	GENERIC(
		SIZE : INTEGER := 32
	);
	PORT ( S 		: IN STD_LOGIC_VECTOR(2 DOWNTO 0) ;
			A, B 		: IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) ;
			F 			: BUFFER STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) ;
			COMPARE	: OUT STD_LOGIC ) ;
END ALU ;

ARCHITECTURE BEHAVIOR OF ALU IS
	BEGIN
	PROCESS ( S, A, B )
	BEGIN
		CASE S IS
			WHEN "000" =>
			F <= x"00000000" ;
			WHEN "001" =>
			F <= B - A ;
			WHEN "010" =>
			F <= A - B ;
			WHEN "011" =>
			F <= A + B ;
			WHEN "100" =>
			F <= A XOR B ;
			WHEN "101" =>
			F <= A OR B ;
			WHEN "110" =>
			F <= A AND B ;
			WHEN OTHERS =>
			F <= x"11111111" ;
			--COMPARE <= '0';
		END CASE ;
	END PROCESS ;

	PROCESS(F,s)
	BEGIN
		IF (F = x"00000000" AND S = "100") THEN
			COMPARE <= '1';
		ELSE
			COMPARE <= '0';
		END IF;
	END PROCESS;
END BEHAVIOR;

