LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY ADDER IS
	GENERIC (
		SIZE : INTEGER := 32
		);
		
	PORT (
		ADDR_IN : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := "00000000000000000000000000000000";
		ADDR_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := "00000000000000000000000000000000");
END ADDER;

ARCHITECTURE RTL OF ADDER IS

BEGIN

	PROC : PROCESS (ADDR_IN) 
	BEGIN
		ADDR_OUT <= ADDR_IN + 1;
	END PROCESS;
END RTL;
