LIBRARY  IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY D_FF IS 
    PORT (CLK : IN STD_LOGIC := '0';
          EN : IN STD_LOGIC := '0';
			 IDLE : IN STD_LOGIC;
          D   : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
			 LOAD : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
          OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000"
    );
END D_FF;

ARCHITECTURE RTL OF D_FF IS
BEGIN
   proc_name: process(CLK,EN)
   begin
       if (RISING_EDGE(CLK)) then
          IF (EN = '1' AND IDLE = '0') THEN  
					OUTPUT <= D;
			 ELSIF (EN = '0' AND IDLE = '1') THEN
					OUTPUT <= LOAD;
			 END IF;
		 END IF;
   end process proc_name;
	
END RTL;




