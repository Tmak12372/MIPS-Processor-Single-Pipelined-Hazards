LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TESTBENCH IS
END TESTBENCH;

ARCHITECTURE RTL OF TESTBENCH IS
COMPONENT MIPS_PROCESSOR IS
	GENERIC(
		SIZE : INTEGER := 32
		);
	PORT (
		CLK 			: IN STD_LOGIC;
		FORA,FORB 	: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		INSTRUCTION : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		ALU_OUT		: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		DATA_OUT    : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		PC    		: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);

END COMPONENT;
	
	
	SIGNAL CLK_TB,STOP_BIT : STD_LOGIC;
	SIGNAL FORA_TB,FORB_TB : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL INSTRUCTION_OUT_TB : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ALU_OUT_TB,DATA_OUT_TB,PC_ADDRESS_TB : STD_LOGIC_VECTOR(6 DOWNTO 0);
BEGIN

	UUT : MIPS_PROCESSOR PORT MAP(CLK_TB,FORA_TB,FORB_TB,INSTRUCTION_OUT_TB,ALU_OUT_TB,DATA_OUT_TB,PC_ADDRESS_TB);

	CLK_1 : PROCESS
		BEGIN
			CLK_TB <= '1'; WAIT FOR 10NS;
			CLK_TB <= '0'; WAIT FOR 10NS;
			IF (STOP_BIT = '1') THEN
				WAIT;
			END IF;
			
	END PROCESS;
	
	STIMULUS : PROCESS
	BEGIN
		WAIT FOR 500NS;
		STOP_BIT <= '1'; --USED FOR GOING THROUGH INSTRUCTIONS
		WAIT;
	END PROCESS;
END RTL;