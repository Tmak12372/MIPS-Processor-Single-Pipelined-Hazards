LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY ADDER IS
	GENERIC (
		SIZE : INTEGER := 32
		);
	PORT (
		ADDRESS_IN  : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := (OTHERS => '0');
		ADDRESS_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := (OTHERS => '0')
		);
END ADDER;

ARCHITECTURE RTL OF ADDER IS
BEGIN
	PROC : PROCESS (ADDRESS_IN) 
	BEGIN
		ADDRESS_OUT <= ADDRESS_IN + 4;  --Increment the Program counter by 1 I chose 1 since my .mif file is incremented address by 1
	END PROCESS;
END RTL;
