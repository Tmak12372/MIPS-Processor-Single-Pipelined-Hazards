LIBRARY  IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY MUX_32_1 IS 
    PORT (
    SEL : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    IN1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN5 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN6 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN7 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN8 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN9 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN13 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN14 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN15 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN16 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN17 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN18 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN19 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN23 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN24 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN25 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN26 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN27 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN28 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN29 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN30 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN31 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN32 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END MUX_32_1;



ARCHITECTURE RTL OF MUX_32_1 IS
BEGIN
    OUTPUT <= IN1 WHEN SEL = "00000"; --1
    OUTPUT <= IN2 WHEN SEL = "00001"; --2
    OUTPUT <= IN3 WHEN SEL = "00010"; --3
    OUTPUT <= IN4 WHEN SEL = "00011"; --4
    OUTPUT <= IN5 WHEN SEL = "00100"; --5
    OUTPUT <= IN6 WHEN SEL = "00101"; --6
    OUTPUT <= IN7 WHEN SEL = "00110"; --7
    OUTPUT <= IN8 WHEN SEL = "00111"; --8
    OUTPUT <= IN9 WHEN SEL = "01000"; --9
    OUTPUT <= IN10 WHEN SEL = "01001"; --10
    OUTPUT <= IN11 WHEN SEL = "01010"; --11
    OUTPUT <= IN12 WHEN SEL = "01011"; --12
    OUTPUT <= IN13 WHEN SEL = "01100"; --13
    OUTPUT <= IN14 WHEN SEL = "01101"; --14
    OUTPUT <= IN15 WHEN SEL = "01110"; --15
    OUTPUT <= IN16 WHEN SEL = "01111"; --16
    OUTPUT <= IN17 WHEN SEL = "10000"; --17
    OUTPUT <= IN18 WHEN SEL = "10001"; --18
    OUTPUT <= IN19 WHEN SEL = "10010"; --19
    OUTPUT <= IN20 WHEN SEL = "10011"; --20
    OUTPUT <= IN21 WHEN SEL = "10100"; --21
    OUTPUT <= IN22 WHEN SEL = "10101"; --22
    OUTPUT <= IN23 WHEN SEL = "10110"; --23
    OUTPUT <= IN24 WHEN SEL = "10111"; --24
    OUTPUT <= IN25 WHEN SEL = "11000"; --25
    OUTPUT <= IN26 WHEN SEL = "11001"; --26
    OUTPUT <= IN27 WHEN SEL = "11010"; --27
    OUTPUT <= IN28 WHEN SEL = "11011"; --28
    OUTPUT <= IN29 WHEN SEL = "11100"; --29
    OUTPUT <= IN30 WHEN SEL = "11101"; --30
    OUTPUT <= IN31 WHEN SEL = "11110"; --31
    OUTPUT <= IN32 WHEN SEL = "11111"; --32
END RTL;

