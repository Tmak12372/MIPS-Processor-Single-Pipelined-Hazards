LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX IS
	GENERIC(
		SIZE : INTEGER := 32
	);
	port(
		SEL			: IN STD_LOGIC;
		INPUT_0		: IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		INPUT_1  	: IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		OUTPUT		: OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)
	);
		
END MUX;


ARCHITECTURE RTL OF MUX IS
BEGIN

	PROCESS (SEL,INPUT_0,INPUT_1)
	BEGIN
		CASE SEL IS
			WHEN '0' => OUTPUT <= INPUT_0;
			WHEN '1' => OUTPUT <= INPUT_1; -- FOR SIGN_EXTENDED
			WHEN OTHERS => OUTPUT <= INPUT_0;
		END CASE;
	END PROCESS;
END RTL;
