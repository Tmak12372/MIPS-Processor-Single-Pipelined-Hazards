LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TESTBENCH IS
END TESTBENCH;

ARCHITECTURE RTL OF TESTBENCH IS
	COMPONENT MIPS_PROCESSOR IS
		GENERIC(
			SIZE : INTEGER := 32
			);
		PORT (
			CLK : IN STD_LOGIC;
			INSTRUCTION_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)
			);

	END COMPONENT;
	
	
	SIGNAL CLK_TB : STD_LOGIC;
	SIGNAL INSTRUCTION_OUT_TB : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
	INSTRUCTION_OUT_TB <= "00000000000000000000000000000000";
	UUT : MIPS_PROCESSOR PORT MAP(CLK_TB,INSTRUCTION_OUT_TB);

	CLK_1 : PROCESS
		BEGIN
			
			CLK_TB <= '1'; WAIT FOR 10NS;
			CLK_TB <= '0'; WAIT FOR 10NS;
	END PROCESS;
	
	STIMULUS : PROCESS
	BEGIN
		
		WAIT FOR 100NS;
		WAIT;
	END PROCESS;
	
END RTL;