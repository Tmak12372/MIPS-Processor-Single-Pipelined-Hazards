LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY MEM_WB IS
	GENERIC(
		SIZE : INTEGER := 32
		);
	PORT (CLK : IN STD_LOGIC;
			RESET : IN STD_LOGIC;
			WB : IN STD_LOGIC_VECTOR(1 DOWNTO 0);	
			READ_DATA : IN  STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			ALU_RESULT : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			MUX_RESULT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			WB_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);	
			READ_DATA_OUT : OUT  STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			ALU_RESULT_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			MUX_RESULT_OUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
			);
END MEM_WB;


ARCHITECTURE RTL OF MEM_WB IS
BEGIN
	PROC : PROCESS(CLK)
	BEGIN
		IF (RISING_EDGE(CLK)) THEN
			IF (RESET = '0') THEN
				WB_OUT <= WB;
				READ_DATA_OUT <= READ_DATA;
				ALU_RESULT_OUT <= ALU_RESULT;
				MUX_RESULT_OUT <= MUX_RESULT;
			ELSE
				WB_OUT <= (OTHERS => '0');
				READ_DATA_OUT <= (OTHERS => '0');
				ALU_RESULT_OUT <= (OTHERS => '0');
				MUX_RESULT_OUT <= (OTHERS => '0');
			END IF;
		END IF;
	END PROCESS;
END RTL;