LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY PROGRAM_COUNTER IS
	GENERIC (
		SIZE : INTEGER := 32
		);
		
	PORT (
		CLK 		: IN STD_LOGIC;
		RES		: IN STD_LOGIC;
		ADDR_IN  : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := "00000000000000000000000000000000";
		ADDR_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := "00000000000000000000000000000000");
END PROGRAM_COUNTER;

ARCHITECTURE RTL OF PROGRAM_COUNTER IS

BEGIN

	PROC : PROCESS (CLK,RES) 
	BEGIN
		IF (RES = '1') THEN
			ADDR_OUT <= "00000000000000000000000000000000";
		ELSIF (RISING_EDGE(CLK)) THEN
				ADDR_OUT <= ADDR_IN;
		END IF;
	END PROCESS;
END RTL;
