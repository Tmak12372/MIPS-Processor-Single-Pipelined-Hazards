LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SIGN_EXTEND IS
	GENERIC(
		SIZE : INTEGER := 32
	);
	port(
		INPUT		: IN STD_LOGIC_VECTOR(SIZE-17 DOWNTO 0);
		OUTPUT	: OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0));
		
END SIGN_EXTEND;

ARCHITECTURE RTL of SIGN_EXTEND IS
	
	BEGIN
	PROCESS(INPUT)
	BEGIN
		CASE INPUT(15) IS
			WHEN '1' => OUTPUT <= ("1111111111111111" & INPUT);
			WHEN '0' => OUTPUT <= ("0000000000000000" & INPUT);
			WHEN OTHERS => OUTPUT <= ("0000000000000000" & INPUT);
		END CASE;
	END PROCESS;
END RTL;