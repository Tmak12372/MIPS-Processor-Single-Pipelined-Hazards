LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TESTBENCH IS
END TESTBENCH;

ARCHITECTURE RTL OF TESTBENCH IS
COMPONENT MIPS_PROCESSOR IS
	GENERIC(
		SIZE : INTEGER := 32
		);
	PORT (
		CLK 		: IN STD_LOGIC;
		REG_WRITE_TO_TB : OUT STD_LOGIC;
		REG_DEST_TO_TB : OUT STD_LOGIC;
		MEMTOREG_TO_TB : OUT STD_LOGIC;
		ALU_SRC_TO_TB : OUT STD_LOGIC;
		ALU_OP_TO_TB : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		MEMREAD_TO_TB : OUT STD_LOGIC;
		MEMWRITE_TO_TB : OUT STD_LOGIC;
		BRANCH_TO_TB  : OUT STD_LOGIC;
		BRANCH_TAKEN : OUT STD_LOGIC;
		ALU_RESULT_TO_TB : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		WRITE_DATA_TO_TB : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		READ_DATA_DM_TO_TB : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		INSTRUCTION : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)
		);

END COMPONENT;
	
	
	SIGNAL CLK_TB,REG_WRITE_TB,ALU_SRC_TB,MEMTOREG_TB,MEMREAD_TB,MEMWRITE_TB,BRANCH_TB,BRANCH_TAKEN_TB,REG_DEST_TB,STOP_BIT : STD_LOGIC;
	SIGNAL ALU_OP_TB : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL INSTRUCTION_TB,READ_DATA_DM_TB,WRITE_DATA_TB,ALU_RESULT_TB : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN

	UUT : MIPS_PROCESSOR PORT MAP(CLK_TB,REG_WRITE_TB,REG_DEST_TB,MEMTOREG_TB,ALU_SRC_TB,ALU_OP_TB,MEMREAD_TB,MEMWRITE_TB,BRANCH_TB,BRANCH_TAKEN_TB,ALU_RESULT_TB,WRITE_DATA_TB,READ_DATA_DM_TB,INSTRUCTION_TB);

	CLK_1 : PROCESS
		BEGIN
			CLK_TB <= '1'; WAIT FOR 10NS;
			CLK_TB <= '0'; WAIT FOR 10NS;
			IF (STOP_BIT = '1') THEN
				WAIT;
			END IF;
			
	END PROCESS;
	
	STIMULUS : PROCESS
	BEGIN
		WAIT FOR 500NS;
		STOP_BIT <= '1'; --USED FOR GOING THROUGH INSTRUCTIONS
		WAIT;
	END PROCESS;
END RTL;