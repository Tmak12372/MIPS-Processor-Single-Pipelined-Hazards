LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALU IS
	GENERIC(
		SIZE : INTEGER := 32
	);
	PORT ( S : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
			A, B : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) ;
			SHIFT_AMOUNT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			F : BUFFER STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) ;
			COMPARE: OUT STD_LOGIC ) ;
END ALU ;

ARCHITECTURE BEHAVIOR OF ALU IS
	BEGIN
	PROCESS ( S, A, B, SHIFT_AMOUNT )
	BEGIN
		CASE S IS
			WHEN "0110" =>
			F <= A - B ;
			WHEN "0010" =>
			F <= A + B ;
			WHEN "0001" =>
			F <= A OR B ;
			WHEN "0000" =>
			F <= A AND B ;
			WHEN "1100" =>
			F <= A NOR B ;
			WHEN "0111" =>
			F <= A XOR B ;
--			WHEN "1010" =>
--				IF (A < B) THEN
--					F <= x"00000001";
--				ELSE
--					F <= x"00000000";
--				END IF;
			WHEN "1011" =>
			F <= STD_LOGIC_VECTOR(unsigned(B) SLL TO_INTEGER(UNSIGNED(SHIFT_AMOUNT)));
--			WHEN "1100" =>
--				F <= STD_LOGIC_VECTOR(unsigned(B) SRL TO_INTEGER(UNSIGNED(SHIFT_AMOUNT)));
			WHEN OTHERS =>
			F <= x"00000000" ;
			--COMPARE <= '0';
		END CASE ;
	END PROCESS ;

	PROCESS(F,s)
	BEGIN
		IF ((F = x"00000000")) THEN
			COMPARE <= '1';
		ELSE
			COMPARE <= '0';
		END IF;
	END PROCESS;
END BEHAVIOR;

