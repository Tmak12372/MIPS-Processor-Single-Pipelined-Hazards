LIBRARY  IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY MUX_32_1 IS 
    PORT (
    SEL : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    IN1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN5 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN6 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN7 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN8 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN9 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN13 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN14 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN15 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN16 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN17 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN18 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN19 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN23 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN24 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN25 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN26 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN27 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN28 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN29 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN30 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN31 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN32 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END MUX_32_1;



ARCHITECTURE RTL OF MUX_32_1 IS
BEGIN
    OUTPUT <= IN1 WHEN SEL = "00000" ELSE
				  IN2 WHEN SEL = "00001" ELSE
				  IN3 WHEN SEL = "00010" ELSE
				  IN4 WHEN SEL = "00011" ELSE
				  IN5 WHEN SEL = "00100" ELSE
				  IN6 WHEN SEL = "00101" ELSE
				  IN7 WHEN SEL = "00110" ELSE
				  IN8 WHEN SEL = "00111" ELSE
				  IN9 WHEN SEL = "01000" ELSE
				  IN10 WHEN SEL = "01001" ELSE
				  IN11 WHEN SEL = "01010" ELSE
				  IN12 WHEN SEL = "01011" ELSE
				  IN13 WHEN SEL = "01100" ELSE
				  IN14 WHEN SEL = "01101" ELSE
				  IN15 WHEN SEL = "01110" ELSE
				  IN16 WHEN SEL = "01111" ELSE
				  IN17 WHEN SEL = "10000" ELSE
				  IN18 WHEN SEL = "10001" ELSE
				  IN19 WHEN SEL = "10010" ELSE
				  IN20 WHEN SEL = "10011" ELSE
				  IN21 WHEN SEL = "10100" ELSE
				  IN22 WHEN SEL = "10101" ELSE
				  IN23 WHEN SEL = "10110" ELSE
				  IN24 WHEN SEL = "10111" ELSE
				  IN25 WHEN SEL = "11000" ELSE
				  IN26 WHEN SEL = "11001" ELSE
				  IN27 WHEN SEL = "11010" ELSE
				  IN28 WHEN SEL = "11011" ELSE
				  IN29 WHEN SEL = "11100" ELSE
				  IN30 WHEN SEL = "11101" ELSE
				  IN31 WHEN SEL = "11110" ELSE
				  IN32 WHEN SEL = "11111" ELSE
				  IN1;
END RTL;

