LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
LIBRARY WORK;

ENTITY REGISTERS IS
	GENERIC(
		SIZE : INTEGER := 32
	);
	PORT(
		CLK																		: IN STD_LOGIC := '0';
		RES																		: IN STD_LOGIC := '0';
		REGWRITE																	: IN STD_LOGIC := '0';
		READ_REGISTER_1, READ_REGISTER_2, WRITE_REGISTER			: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		WRITE_DATA																: IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0) := "00000000000000000000000000000000";
		READ_DATA_1, READ_DATA_2											: OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)
	);
END REGISTERS;

ARCHITECTURE RTL OF REGISTERS IS
COMPONENT Decoder_5_32 IS 
    PORT (INPUT : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
          OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END COMPONENT;

COMPONENT D_FF IS 
    PORT (CLK : IN STD_LOGIC := '0';
          EN : IN STD_LOGIC := '0';
			 IDLE : IN STD_LOGIC;
          D   : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
			 LOAD : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
          OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000"
    );
END COMPONENT;

COMPONENT MUX_32_1 IS 
    PORT (
    SEL : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    IN1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN5 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN6 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN7 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN8 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN9 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN13 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN14 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN15 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN16 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN17 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN18 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN19 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN23 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN24 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN25 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN26 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN27 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN28 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN29 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN30 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN31 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IN32 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END COMPONENT;


COMPONENT REGISTER_AND IS 
    PORT (A : IN STD_LOGIC;
          B   : IN STD_LOGIC;
          F : OUT STD_LOGIC
    );
END COMPONENT;

SIGNAL DECODER_OUTPUT : STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";


TYPE MATRIX IS ARRAY(0 TO SIZE-1) OF STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
	SIGNAL Registers : MATRIX := (OTHERS => (OTHERS => '0'));								 

TYPE MATRIX1 IS ARRAY(0 TO SIZE-1) OF STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
	SIGNAL Registers1 : MATRIX := (OTHERS => (OTHERS => '0'));
								 
								 
								 
								 
TYPE MAT IS ARRAY(0 TO SIZE-1) OF STD_LOGIC;
	SIGNAL C : MAT := (OTHERS => '0');
								





	signal IsStartup : STD_LOGIC := '1';

BEGIN
	
	process(CLK,RES)
	begin
	  if (rising_edge(CLK)) then
		  IF RES = '0' THEN
				IsStartup <= '0';
		  else 
				IsStartup <= '1';
		  END IF;
	  end if;  
	end process;
	
	
    U50 : Decoder_5_32 PORT MAP (WRITE_REGISTER,DECODER_OUTPUT);

	 GEN1 : for i in 0 to 31 generate
		U51 : REGISTER_AND PORT MAP(REGWRITE,DECODER_OUTPUT(i),C(i));
	 end generate;
	 
	 GEN2 : for i in 0 to 31 generate
		U90 : D_FF PORT MAP (CLK,C(i),IsStartup,WRITE_DATA,REGISTERS1(i),REGISTERS(i));
	 end generate;
	 
    U122 : MUX_32_1 PORT MAP (READ_REGISTER_1,REGISTERS(0),REGISTERS(1),REGISTERS(2),REGISTERS(3),REGISTERS(4),REGISTERS(5),REGISTERS(6),REGISTERS(7),REGISTERS(8),REGISTERS(9),REGISTERS(10),REGISTERS(11),REGISTERS(12),REGISTERS(13),REGISTERS(14),REGISTERS(15),REGISTERS(16),REGISTERS(17),REGISTERS(18),REGISTERS(19),REGISTERS(20),REGISTERS(21),REGISTERS(22),REGISTERS(23),REGISTERS(24),REGISTERS(25),REGISTERS(26),REGISTERS(27),REGISTERS(28),REGISTERS(29),REGISTERS(30),REGISTERS(31),READ_DATA_1);
    U123 : MUX_32_1 PORT MAP (READ_REGISTER_2,REGISTERS(0),REGISTERS(1),REGISTERS(2),REGISTERS(3),REGISTERS(4),REGISTERS(5),REGISTERS(6),REGISTERS(7),REGISTERS(8),REGISTERS(9),REGISTERS(10),REGISTERS(11),REGISTERS(12),REGISTERS(13),REGISTERS(14),REGISTERS(15),REGISTERS(16),REGISTERS(17),REGISTERS(18),REGISTERS(19),REGISTERS(20),REGISTERS(21),REGISTERS(22),REGISTERS(23),REGISTERS(24),REGISTERS(25),REGISTERS(26),REGISTERS(27),REGISTERS(28),REGISTERS(29),REGISTERS(30),REGISTERS(31),READ_DATA_2);
	 
	 
	 
	 END RTL;