LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY ID_EX IS
	GENERIC(
		SIZE : INTEGER := 32
		);
	PORT (CLK : IN STD_LOGIC;
			RESET : IN STD_LOGIC;
			BNE : IN STD_LOGIC;
			WB : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			M : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			EX : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			PC : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			READ_DATA_1_IN : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			READ_DATA_2_IN : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			SIGN_EXTEND : IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			INST2016 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			INST1511 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			WB_OUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
			M_OUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
			EX_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			PC_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			READ_DATA_1_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			READ_DATA_2_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			SIGN_EXTEND_OUT : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
			INST2016_OUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			INST1511_OUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			BNE_OUT : OUT STD_LOGIC
			);
END ID_EX;

ARCHITECTURE RTL OF ID_EX IS
BEGIN
	PROC : PROCESS(CLK)
	BEGIN
		IF (RISING_EDGE(CLK)) THEN
			IF (RESET = '0') THEN
				WB_OUT <= WB;
				M_OUT <= M;
				EX_OUT <= EX;
				PC_OUT <= PC;
				READ_DATA_1_OUT <= READ_DATA_1_IN;
				READ_DATA_2_OUT <= READ_DATA_2_IN;
				SIGN_EXTEND_OUT <= SIGN_EXTEND;
				INST2016_OUT <= INST2016;
				INST1511_OUT <= INST1511;
				BNE_OUT <= BNE;
			ELSE
				WB_OUT <= (OTHERS => '0');
				M_OUT <= (OTHERS => '0');
				EX_OUT <= (OTHERS => '0');
				PC_OUT <= (OTHERS => '0');
				READ_DATA_1_OUT <= (OTHERS => '0');
				READ_DATA_2_OUT <= (OTHERS => '0');
				SIGN_EXTEND_OUT <= (OTHERS => '0');
				INST2016_OUT <= (OTHERS => '0');
				INST1511_OUT <= (OTHERS => '0');
				BNE_OUT <= '0';
			END IF;
		END IF;
	END PROCESS;
END RTL;
	
	