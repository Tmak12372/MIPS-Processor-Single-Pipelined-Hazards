LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
LIBRARY WORK;

ENTITY REGISTERS IS
	GENERIC(
		SIZE : INTEGER := 32
	);
	PORT(
		CLK																		: IN STD_LOGIC;
		REGWRITE																	: IN STD_LOGIC;
		READ_REGISTER_1, READ_REGISTER_2, WRITE_REGISTER			: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		WRITE_DATA																: IN STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		READ_DATA_1, READ_DATA_2											: OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0)
	);
END REGISTERS;

ARCHITECTURE RTL OF REGISTERS IS
SIGNAL DECODER_OUTPUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG1_CLK : STD_LOGIC;
SIGNAL REG2_CLK : STD_LOGIC;
SIGNAL REG3_CLK : STD_LOGIC;
SIGNAL REG4_CLK : STD_LOGIC;
SIGNAL REG5_CLK : STD_LOGIC;
SIGNAL REG6_CLK : STD_LOGIC;
SIGNAL REG7_CLK : STD_LOGIC;
SIGNAL REG8_CLK : STD_LOGIC;
SIGNAL REG9_CLK : STD_LOGIC;
SIGNAL REG10_CLK : STD_LOGIC;
SIGNAL REG11_CLK : STD_LOGIC;
SIGNAL REG12_CLK : STD_LOGIC;
SIGNAL REG13_CLK : STD_LOGIC;
SIGNAL REG14_CLK : STD_LOGIC;
SIGNAL REG15_CLK : STD_LOGIC;
SIGNAL REG16_CLK : STD_LOGIC;
SIGNAL REG17_CLK : STD_LOGIC;
SIGNAL REG18_CLK : STD_LOGIC;
SIGNAL REG19_CLK : STD_LOGIC;
SIGNAL REG20_CLK : STD_LOGIC;
SIGNAL REG21_CLK : STD_LOGIC;
SIGNAL REG22_CLK : STD_LOGIC;
SIGNAL REG23_CLK : STD_LOGIC;
SIGNAL REG24_CLK : STD_LOGIC;
SIGNAL REG25_CLK : STD_LOGIC;
SIGNAL REG26_CLK : STD_LOGIC;
SIGNAL REG27_CLK : STD_LOGIC;
SIGNAL REG28_CLK : STD_LOGIC;
SIGNAL REG29_CLK : STD_LOGIC;
SIGNAL REG30_CLK : STD_LOGIC;
SIGNAL REG31_CLK : STD_LOGIC;
SIGNAL REG32_CLK : STD_LOGIC;
SIGNAL REG1_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG2_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG3_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG4_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG5_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG6_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG7_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG8_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG9_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG10_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG11_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG12_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG13_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG14_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG15_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG16_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG17_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG18_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG19_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG20_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG21_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG22_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG23_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG24_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG25_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG26_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG27_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG28_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG29_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG30_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG31_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG32_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
    U50 : WORK.Decoder_5_32 PORT MAP (WRITE_REGISTER,DECODER_OUTPUT);

    U51 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(0),REG1_CLK);
    U52 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(1),REG2_CLK);
    U53 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(2),REG3_CLK);
    U54 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(3),REG4_CLK);
    U55 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(4),REG5_CLK);
    U56 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(5),REG6_CLK);
    U57 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(6),REG7_CLK);
    U58 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(7),REG8_CLK);
    U59 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(8),REG9_CLK);
    U60 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(9),REG10_CLK);
    U61 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(10),REG11_CLK);
    U62 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(11),REG12_CLK);
    U63 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(12),REG13_CLK);
    U64 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(13),REG14_CLK);
    U65 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(14),REG15_CLK);
    U66 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(15),REG16_CLK);
    U67 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(16),REG17_CLK);
    U68 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(17),REG18_CLK);
    U69 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(18),REG19_CLK);
    U70 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(19),REG20_CLK);
    U71 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(20),REG21_CLK);
    U72 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(21),REG22_CLK);
    U73 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(22),REG23_CLK);
    U74 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(23),REG24_CLK);
    U75 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(24),REG25_CLK);
    U76 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(25),REG26_CLK);
    U77 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(26),REG27_CLK);
    U78 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(27),REG28_CLK);
    U79 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(28),REG29_CLK);
    U80 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(29),REG30_CLK);
    U81 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(30),REG31_CLK);
    U82 : WORK.REGISTER_AND PORT MAP (WRITE_DATA,DECODER_OUTPUT(31),REG32_CLK);

    U90 : WORK.D_FF PORT MAP (CLK,REG1_CLK,WRITE_DATA,REG1_VALUE);
    U91 : WORK.D_FF PORT MAP (CLK,REG2_CLK,WRITE_DATA,REG2_VALUE);
    U92 : WORK.D_FF PORT MAP (CLK,REG3_CLK,WRITE_DATA,REG3_VALUE);
    U93 : WORK.D_FF PORT MAP (CLK,REG4_CLK,WRITE_DATA,REG4_VALUE);
    U94 : WORK.D_FF PORT MAP (CLK,REG5_CLK,WRITE_DATA,REG5_VALUE);
    U95 : WORK.D_FF PORT MAP (CLK,REG6_CLK,WRITE_DATA,REG6_VALUE);
    U96 : WORK.D_FF PORT MAP (CLK,REG7_CLK,WRITE_DATA,REG7_VALUE);
    U97 : WORK.D_FF PORT MAP (CLK,REG8_CLK,WRITE_DATA,REG8_VALUE);
    U98 : WORK.D_FF PORT MAP (CLK,REG9_CLK,WRITE_DATA,REG9_VALUE);
    U99 : WORK.D_FF PORT MAP (CLK,REG10_CLK,WRITE_DATA,REG10_VALUE);
    U100 : WORK.D_FF PORT MAP (CLK,REG11_CLK,WRITE_DATA,REG11_VALUE);
    U101 : WORK.D_FF PORT MAP (CLK,REG12_CLK,WRITE_DATA,REG12_VALUE);
    U102 : WORK.D_FF PORT MAP (CLK,REG13_CLK,WRITE_DATA,REG13_VALUE);
    U103 : WORK.D_FF PORT MAP (CLK,REG14_CLK,WRITE_DATA,REG14_VALUE);
    U104 : WORK.D_FF PORT MAP (CLK,REG15_CLK,WRITE_DATA,REG15_VALUE);
    U105 : WORK.D_FF PORT MAP (CLK,REG16_CLK,WRITE_DATA,REG16_VALUE);
    U106 : WORK.D_FF PORT MAP (CLK,REG17_CLK,WRITE_DATA,REG17_VALUE);
    U107 : WORK.D_FF PORT MAP (CLK,REG18_CLK,WRITE_DATA,REG18_VALUE);
    U108 : WORK.D_FF PORT MAP (CLK,REG19_CLK,WRITE_DATA,REG19_VALUE);
    U109 : WORK.D_FF PORT MAP (CLK,REG20_CLK,WRITE_DATA,REG20_VALUE);
    U110 : WORK.D_FF PORT MAP (CLK,REG21_CLK,WRITE_DATA,REG21_VALUE);
    U111 : WORK.D_FF PORT MAP (CLK,REG22_CLK,WRITE_DATA,REG22_VALUE);
    U112 : WORK.D_FF PORT MAP (CLK,REG23_CLK,WRITE_DATA,REG23_VALUE);
    U113 : WORK.D_FF PORT MAP (CLK,REG24_CLK,WRITE_DATA,REG24_VALUE);
    U114 : WORK.D_FF PORT MAP (CLK,REG25_CLK,WRITE_DATA,REG25_VALUE);
    U115 : WORK.D_FF PORT MAP (CLK,REG26_CLK,WRITE_DATA,REG26_VALUE);
    U116 : WORK.D_FF PORT MAP (CLK,REG27_CLK,WRITE_DATA,REG27_VALUE);
    U117 : WORK.D_FF PORT MAP (CLK,REG28_CLK,WRITE_DATA,REG28_VALUE);
    U118 : WORK.D_FF PORT MAP (CLK,REG29_CLK,WRITE_DATA,REG29_VALUE);
    U119 : WORK.D_FF PORT MAP (CLK,REG30_CLK,WRITE_DATA,REG30_VALUE);
    U120 : WORK.D_FF PORT MAP (CLK,REG31_CLK,WRITE_DATA,REG31_VALUE);
    U121 : WORK.D_FF PORT MAP (CLK,REG32_CLK,WRITE_DATA,REG32_VALUE);

    U122 : WORK.MUX_32_1 PORT MAP (READ_REGISTER_1,REG1_VALUE,REG2_VALUE,REG3_VALUE,REG4_VALUE,REG5_VALUE,REG6_VALUE,REG7_VALUE,REG8_VALUE,REG9_VALUE,REG10_VALUE,REG11_VALUE,REG12_VALUE,REG13_VALUE,REG14_VALUE,REG15_VALUE,REG16_VALUE,REG17_VALUE,REG18_VALUE,REG19_VALUE,REG20_VALUE,REG21_VALUE,REG22_VALUE,REG23_VALUE,REG24_VALUE,REG25_VALUE,REG26_VALUE,REG27_VALUE,REG28_VALUE,REG29_VALUE,REG30_VALUE,REG31_VALUE,REG32_VALUE,READ_DATA_1);
    U123 : WORK.MUX_32_1 PORT MAP (READ_REGISTER_2,REG1_VALUE,REG2_VALUE,REG3_VALUE,REG4_VALUE,REG5_VALUE,REG6_VALUE,REG7_VALUE,REG8_VALUE,REG9_VALUE,REG10_VALUE,REG11_VALUE,REG12_VALUE,REG13_VALUE,REG14_VALUE,REG15_VALUE,REG16_VALUE,REG17_VALUE,REG18_VALUE,REG19_VALUE,REG20_VALUE,REG21_VALUE,REG22_VALUE,REG23_VALUE,REG24_VALUE,REG25_VALUE,REG26_VALUE,REG27_VALUE,REG28_VALUE,REG29_VALUE,REG30_VALUE,REG31_VALUE,REG32_VALUE,READ_DATA_2);