LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TESTBENCH IS
END TESTBENCH;

ARCHITECTURE RTL OF TESTBENCH IS
COMPONENT MIPS_PROCESSOR IS
	GENERIC(
		SIZE : INTEGER := 32
		);
	PORT (
		CLK 		: IN STD_LOGIC;
--		SEL		: IN STD_LOGIC;
		INSTRUCTION : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		ALU_RES   : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		DATA1,DATA2   : OUT STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);
		CONTROL : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
--		dFix         : OUT STD_LOGIC_VECTOR(5 downto 0) := "111111";
--		ledFix       : OUT STD_LOGIC_VECTOR(9 downto 0) := "0000000000";
--		hex5         : OUT STD_LOGIC_VECTOR(6 downto 0);
--		hex4         : OUT STD_LOGIC_VECTOR(6 downto 0);
--		hex3         : OUT STD_LOGIC_VECTOR(6 downto 0);
--		hex2         : OUT STD_LOGIC_VECTOR(6 downto 0);
--		hex1         : OUT STD_LOGIC_VECTOR(6 downto 0);
--		hex0         : OUT STD_LOGIC_VECTOR(6 downto 0)
		);

END COMPONENT;
	
	
	SIGNAL CLK_TB,STOP_BIT : STD_LOGIC;
	SIGNAL CONTROL_TB : STD_LOGIC_VECTOR(8 DOWNTO 0);
	SIGNAL ALU_RES_TB,INSTRUCTION_TB,DATA1_TB,DATA2_TB : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
	UUT : MIPS_PROCESSOR PORT MAP(CLK_TB,INSTRUCTION_TB,ALU_RES_TB,DATA1_TB,DATA2_TB,CONTROL_TB);

	CLK_1 : PROCESS
		BEGIN
			CLK_TB <= '1'; WAIT FOR 10NS;
			CLK_TB <= '0'; WAIT FOR 10NS;
			IF (STOP_BIT = '1') THEN
				WAIT;
			END IF;
			
	END PROCESS;
	
	STIMULUS : PROCESS
	BEGIN
		
		WAIT FOR 250NS;
		STOP_BIT <= '1'; --USED FOR GOING THROUGH INSTRUCTIONS
		WAIT;
	END PROCESS;
END RTL;