LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY INSTRUCTION_REGISTER IS
	
	GENERIC(
		SIZE : INTEGER := 32
		);
	
	PORT(
		CLK					:	IN STD_LOGIC;
		ADDR_IN			   :	IN STD_LOGIC_Vector(SIZE-1 DOWNTO 0);
		DATA_IN				:	IN STD_LOGIC_Vector(SIZE-1 DOWNTO 0);
		ADDR_OUT			   :	OUT STD_LOGIC_Vector(7 DOWNTO 0);
		INST_OUT 	      :	OUT STD_LOGIC_Vector(SIZE-1 DOWNTO 0)
		);
		
END INSTRUCTION_REGISTER;

ARCHITECTURE RTL OF INSTRUCTION_REGISTER IS
	
	BEGIN
	PROC : PROCESS (CLK)
	BEGIN
		if (CLK'EVENT AND CLK = '1') THEN
			ADDR_OUT <= ADDR_IN(7 DOWNTO 0);
			INST_OUT <= DATA_IN;
		END IF;
		
	END PROCESS;
	
END RTL;