LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY HAZARD_MUX IS
	GENERIC (
		SIZE : INTEGER := 32
	);
	PORT (
		SEL : IN STD_LOGIC;
		REG_WRITE : IN STD_LOGIC;
		MEMTOREG : IN STD_LOGIC;
		BRANCH : IN STD_LOGIC;
		MEMREAD : IN STD_LOGIC;
		MEMWRITE : IN STD_LOGIC;
		REG_DEST : IN STD_LOGIC;
		ALU_OP : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		ALU_SRC : IN STD_LOGIC;
		WB_IN_IDEX : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		M_IDEX : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		EX_IDEX : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END HAZARD_MUX;

ARCHITECTURE RTL OF HAZARD_MUX IS
BEGIN
    PROC : PROCESS (SEL,REG_WRITE,MEMTOREG,BRANCH,MEMREAD,MEMWRITE,REG_DEST,ALU_OP,ALU_SRC) 
	BEGIN
        IF (SEL = '0') THEN
				WB_IN_IDEX(1) <= REG_WRITE;
				WB_IN_IDEX(0) <= MEMTOREG;
				M_IDEX(2) <= BRANCH;
				M_IDEX(1) <= MEMREAD;
				M_IDEX(0) <= MEMWRITE;
				EX_IDEX(3) <= REG_DEST;
				EX_IDEX(2) <= ALU_OP(1);
				EX_IDEX(1) <= ALU_OP(0);
				EX_IDEX(0) <= ALU_SRC;
        ELSE
				WB_IN_IDEX <= "00";
				M_IDEX <= "000";
				EX_IDEX <= "0000";
		  END IF;
    END PROCESS;
END RTL;