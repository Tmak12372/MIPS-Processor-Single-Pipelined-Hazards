LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY HAZARD_UNIT IS
	GENERIC (
		SIZE : INTEGER := 32
	);
	PORT (
        ID_EX_REGISTER_RS  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        ID_EX_REGISTER_RT  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        IF_ID_REGISTER_RS  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        IF_ID_REGISTER_RT  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        ID_EX_MEMREAD      : IN STD_LOGIC;
        PC_WRITE    : OUT STD_LOGIC;
        IF_ID_WRITE : OUT STD_LOGIC;
        MUX_SEL     : OUT STD_LOGIC
    );
END HAZARD_UNIT;

ARCHITECTURE RTL OF HAZARD_UNIT IS
BEGIN
    PROC : PROCESS (ID_EX_REGISTER_RS,ID_EX_REGISTER_RT,ID_EX_MEMREAD) 
	BEGIN
        IF (ID_EX_MEMREAD = '1' AND (ID_EX_REGISTER_RT /= "00000") AND ((ID_EX_REGISTER_RT = IF_ID_REGISTER_RS) OR (ID_EX_REGISTER_RT = IF_ID_REGISTER_RT))) THEN
            PC_WRITE <= '1';
            IF_ID_WRITE <= '1';
            MUX_SEL <= '1';
        ELSE
            PC_WRITE <= '0';
            IF_ID_WRITE <= '0';
            MUX_SEL <= '0';
			END IF;
    END PROCESS;
END RTL;
